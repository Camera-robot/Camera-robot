// This testbench used an image stored in array and produce a VGA stream

`include "img_utils.svh"

module tbench ();

bit reset     = 1'b0;


bit         vga_clk   = 1'b0;// Pixel clock set as 25Mhz
bit         vga_clk2x = 1'b0;// 50Mhz for GeneSync block
logic [9:0] vga_x;         // X position of pixel
logic [8:0] vga_y;         // Y position of pixel
logic       vga_hsync;     // Horizontal Synchro (before every line)
logic       vga_vsync;     // Vertical Synchro (New image on screen)
logic       vga_img;       // img permet de couper r/g/b quand on est hors de l'ecran (back and front porch)

logic [9:0] cam_x;         // X position of pixel in camera
logic [8:0] cam_y;         // Y position of pixel in camera
logic r     ;
logic g     ;
logic b     ;
logic r_out ;
logic g_out ;
logic b_out ;

logic [8:0] X_top;         // X position
logic [8:0] Y_top;         // Y position

// VGA screen is 640x480
// Image Array
pixel_t img_camera [int][int]; // Camera Output is 512x512
pixel_t img_out; // Pixel output after processing
pixel_t img_barycentre;
pixel_t img_vga    [int][int]; // VGA screen is 640x480
pixel_t img_vga_2    [int][int]; // VGA screen is 640x480

// Initialise all array to black
initial begin
  for (int y=0; y < 480; y++) begin
    for (int x=0; x < 640; x++) begin
      img_vga[x][y].b = "00";
      img_vga[x][y].g = "00";
      img_vga[x][y].r = "00";
      img_vga_2[x][y].b = "00";
      img_vga_2[x][y].g = "00";
      img_vga_2[x][y].r = "00";
    end
  end
end

// Le composant vga_sync est un bloc qui g�n�re les signaux HSYNC et VSYNC conform�ment �
// la norme VGA (pour une r�solution de 640x480 pixels). Le signal IMG est � 1 uniquement
// lorsque le canon � �lectrons est dans une zone visible de l'image. Si IMG est � 0, alors
// les signaux R, G et B doivent obligatoirement �tre � 0 aussi. Les signaux X et Y d�signent
// les coordonn�es du pixel de couleurs R, G et B � l'instant consid�r�.
/*vga_sync u_vga_sync (
  .clk   (vga_clk),     // VGA clock (must be set at 25Mhz)
  .rst_n (reset),       // Active Low Reset
  .hsync (vga_hsync),   // VGA Horizontal Synchronisation
  .vsync (vga_vsync),   // VGA Vertical Synchronisation
  .pos_x (vga_x),       // X position of on pixel in the vga screen
  .pos_y (vga_y),       // Y position of on pixel in the vga screen
  .img   (vga_img)      // High when we are inside VGA scree (not in porch of sync area)
);
assign cam_x   = (vga_x > 128 && vga_x < 640) ?  vga_x - 128 : 0; // 128 = 640 (vga) - 512 (camera)
assign cam_y   =                                 vga_y;           // same Y as 512 (canera)  > 480 (vga)
assign cam_img = (vga_x > 128) && vga_img;         // Force vga pixel out of camera to 0*/

/*gensync u_gsync (
  .CLK          (vga_clk),
  .reset        (reset),
  .HSYNC        (vga_hsync),
  .VSYNC        (vga_vsync),
  .IMG          (vga_img),
  .IMGY_out     (),
  .X            (cam_x),
  .Y            (cam_y)
);*/
assign vga_x   = (cam_x < 640) ? cam_x + 128: 0;
assign vga_y   = cam_y;
assign cam_img = vga_img;


top_bar top (
	.CLK_top (vga_clk),
	.reset_top (reset),
	.SW1_top (1'b1),
	.r_top (img_camera[cam_x][cam_y].r), // Input Red Pixel
	.g_top (img_camera[cam_x][cam_y].g), // Input Green Pixel
	.b_top (img_camera[cam_x][cam_y].b), // Input Blue Pixel

	.rout_top (img_barycentre.r),
	.gout_top (img_barycentre.g),
	.bout_top (img_barycentre.b),

	.r_out_proc (img_out.r),
	.g_out_proc (img_out.g),
	.b_out_proc (img_out.b),

	.X_barycentre_top(X_top),
	.Y_barycentre_top(Y_top),

	.HSYNC_top (vga_hsync),
	.VSYNC_top (vga_vsync),
	.cam_x (cam_x),
	.cam_y (cam_y),
	.IMG_top (vga_img)

);



always @(posedge vga_clk) 
  //if ((vga_x < 640) && (vga_y < 480))
  begin
    img_vga[vga_x][vga_y].r = img_out.r & {8{cam_img}};
    img_vga[vga_x][vga_y].g = img_out.g & {8{cam_img}};
    img_vga[vga_x][vga_y].b = img_out.b & {8{cam_img}};

    img_vga_2[vga_x][vga_y].r = img_barycentre.r & {8{cam_img}}; 
    img_vga_2[vga_x][vga_y].g = img_barycentre.g & {8{cam_img}};
    img_vga_2[vga_x][vga_y].b = img_barycentre.b & {8{cam_img}}; 
  end

initial begin
  #103  reset      = 1'b1;
end

// Set Pixel Clock @ 25Mhz --> 40ns
always #20 vga_clk   <= ~vga_clk;
always #10 vga_clk2x <= ~vga_clk2x;

// Read Image From File
initial begin
  read_bmp(img_camera,"/tp/xph3app/xph3app602/Camera_robot/Bench/img/test_bnw_512x512.bmp");//selection image
end

// Write image
initial begin
  @(posedge reset);
  @(posedge vga_vsync);
  @(negedge vga_vsync); 
	write_bmp(img_vga,"img_out.bmp"); // used for detection
  @(posedge vga_vsync);
  @(negedge vga_vsync);
 	write_bmp(img_vga_2,"img_barycentre.bmp"); // used for detection
  @(posedge vga_vsync); 
  @(negedge vga_vsync);
 	write_bmp(img_vga_2,"img_barycentre2.bmp"); // used for detection
  @(posedge vga_vsync); $finish;
end

endmodule
