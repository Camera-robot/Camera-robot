library IEEE;		--à nettoyer en test unitaire à la fin
        use IEEE.std_logic_1164.all;
        use IEEE.std_logic_textio.all;
        use IEEE.std_logic_arith.all;
        use IEEE.numeric_bit.all;
        use IEEE.numeric_std.all;
        use IEEE.std_logic_signed.all;
        use IEEE.std_logic_unsigned.all;
        use IEEE.math_real.all;
        use IEEE.math_complex.all;

library STD;
        use STD.textio;

entity trame_assembler is
	port(	trame_in	:	in	STD_LOGIC_VECTOR(39 downto 0);		--trame avec len + instru + adresse + mvt
		id		:	in	STD_LOGIC_VECTOR(7 downto 0);
		cs		:	in	STD_LOGIC_VECTOR(7 downto 0);
		trame_out	:	out	STD_LOGIC_VECTOR(71 downto 0));
end trame_assembler;

architecture TA of trame_assembler is

	signal header : STD_LOGIC_VECTOR(15 downto 0) := "1111111111111111";

begin
	trame_out <= header & id & trame_in & cs;

end TA;
